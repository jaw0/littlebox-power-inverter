gpi1 output filter


* R @ 56k
* 38V @ 300k


* http://ngspice.sourceforge.net/docs/ngspice23-manual.pdf
*
* 1 3 5
* 2 4 0
*
*
*
*  --+ 1 +--+--+ 3 +--+--
*      L    |    L    |
*                     |
*                     C6
*                     |
*      L    |    L    |
*  --+ 2 +--+--+ 4 +--+--
*

L1 1 3 10u

L2 2 4 10u

L3 3 5 10u

L4 4 0 10u

C6 5 0 .2u

Rload 5 0 1000
Vin   1 2 AC 1000

.AC DEC 1000 10k 10Meg

.control
run
set color0=#fffff0
set color1=black
set color2=#C00000
plot mag(V(5)) loglog
* plot mag(V(5)) loglog xlimit 250k 450k

.endc

.end
