gpi1 output filter

* this is what is on the filter3 board
*
* R @ 14k;  3V @ 300k
*
* 1 3
* 2 0
*
*
*
*  --+ 1 +---+--
*      L     |
*            |
*            C1
*            |
*      L     |
*  --+ 2 +---+--
*


L1 1 3 100u

L2 2 0 100u

C1 3 0 .68u

Rload 3 0 1000
Vin   1 2 AC 1000

.AC DEC 1000 10k 10Meg

.control
run
set color0=#fffff0
set color1=black
set color2=#C00000

plot mag(V(3)) loglog
* plot mag(V(3)) loglog xlimit 250k 650k
.endc

.end
