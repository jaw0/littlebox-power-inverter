gpi1 output filter

* low-pass + notch
* R @ 52k, 157k, 450k, 525k
* ok 290k - 390k; meh @ 600k

* QQQ - use C1+C3; C1+C2; C3+C4 is there a difference?

* http://ngspice.sourceforge.net/docs/ngspice23-manual.pdf
*
* 1 3 5
* 2 4 0
*
*
*      C         C
*  --+ 1 +--+--+ 3 +--+--
*      L    |    L    |
*           |         |
*           C5        C6
*           |         |
*      L    |    L    |
*  --+ 2 +--+--+ 4 +--+--
*                C

L1 1 3 10u
C1 1 3 .027u

L2 2 4 10u

L3 3 5 10u
C3 3 5 .018u

L4 4 0 10u
C4 4 0 .010u

C5 3 4 .1u
C6 5 0 .2u

Rload 5 0 1000
Vin   1 2 AC 1000

.AC DEC 1000 10k 10Meg

.control
run
set color0=#fffff0
set color1=black
set color2=#C00000
plot mag(V(5)) loglog
* plot mag(V(5)) loglog xlimit 250k 450k

.endc

.end
